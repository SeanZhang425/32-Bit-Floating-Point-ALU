/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_ALU (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    wire [7:0] alu_io_out;
    wire [7:0] alu_io_oe;
    
    alu_top u_alu (
        .clk    (clk),
        .rst_n  (rst_n),
        .in     (ui_in),
        .out    (uo_out),
        .io_in  (uio_in),
        .io_out (alu_io_out),
        .io_oe  (alu_io_oe)
    );
        
    assign uio_out = alu_io_out;
    assign uio_oe  = alu_io_oe;
    
    // List all unused inputs to prevent warnings
    wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule
